`ifndef MAC_BW
    `define MAC_BW 12
`endif

`ifndef ACC_DEP
    `define ACC_DEP 4
`endif