`ifndef MAC_BW
    `define MAC_BW 16
`endif