`ifndef MAC_BW
    `define MAC_BW 12
`endif