`ifndef MAC_BW
    `define MAC_BW 20
`endif