`ifndef MAC_BW
    `define MAC_BW 8
`endif